Reverse Breakdown

.include 1N914.txt
.include 1N34A.txt

.option temp = val
Vs 1 0 dc 20
R1 1 2 100
R2 2 0 1k
D1 2 3 1N914
*D1 2 3 1N34A
Vdummy 3 4 dc 0
R3 4 0 100

.dc Vs 0.01 10 0.01 val 20 80 10
.control
run

plot i(Vdummy) vs v(2,3)
meas dc turnon find v(2,3) when i(Vdummy)=1m
meas dc rev_breakdown find v(2,3) when i(Vdummy)=-500u

.endc
.end
