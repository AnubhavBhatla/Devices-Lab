*NMOS Subthreshold slope

.include 2n7000.txt

vgg 1 0 dc 0v
vdd 2 0 dc 5v
vbb 3 0 dc -1.5v
m1 2 1 0 3 2N7000

.dc vgg 0 2 0.01 vbb 0 -1.5 -0.5
.control
run

plot log(-i(vdd))

.endc
.end
