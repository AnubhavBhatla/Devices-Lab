RF Switch Circuit

.include rn142.txt

Vin in 0 sin(0 6 10Meg 0 0)
C1 in 1 100n
R1 1 0 500
D dummy1 1 DRN142S
Vdummy1 2 dummy1 dc 0 ac 0
R2 2 3 500
Vbias 3 0 dc 5
C2 2 out 100n
R3 out dummy2 50
Vdummy2 0 dummy2 dc 0 ac 0

.tran 0.1n 1u
.control
run

plot v(out) v(in)
plot i(Vdummy1) i(Vdummy2)

.endc
.end
