Diode I-V Characteristics

.include rn142.txt

Vs 1 0 dc 20
D1 1 2 DRN142S

R1 2 12 100

V1 12 0 dc 0

.dc Vs 0.01 5 0.01
.control
run

set color0 = white
set color1 = black
set color2 = red

plot i(V1) vs v(1,2)

set color0 = white
set color1 = black
set color2 = red

meas dc cutin find v(1,2) when i(V1) = 1m

plot ln(i(V1)) vs v(1,2)

let derivout = deriv((ln(i(V1))))
meas dc slope find derivout when v(1,2) = 500m

.endc
.end
